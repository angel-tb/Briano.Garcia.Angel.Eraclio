** Profile: "SCHEMATIC1-Amp-Op- no inverso"  [ E:\PRACTICA SCR-TRIAC\Practica-PSpiceFiles\SCHEMATIC1\Amp-Op- no inverso.sim ] 

** Creating circuit file "Amp-Op- no inverso.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 50u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
